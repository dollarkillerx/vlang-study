module main

fn main() {
	nums := [1,2,3]
	println(1 in nums) // in 判断是否包含

	// if p
}