module main

fn main() {
	println("Hello Vlang")
}