module modelt

pub fn add(a int,b int) int {
	return a + b
}