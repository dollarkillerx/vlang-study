module main

fn main() {
	age := 16
	println('you age: $age')

	s := r'hello \n you '  // r 原始字符串
	println('$s')
}