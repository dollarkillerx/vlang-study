module main

fn main() {
	name := 'Bob'
	mut age := 20
	println(name)
	println(age)

	age = 16
	println(age)

	// 默认生成的三常量  加上mut才是常量
}